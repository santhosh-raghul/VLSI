magic
tech scmos
timestamp 1597250001
<< nwell >>
rect -27 -1 29 10
<< polysilicon >>
rect -14 8 -10 12
rect -2 8 2 12
rect 10 8 14 12
rect -14 -29 -10 1
rect -2 -29 2 1
rect 10 -29 14 1
rect -14 -38 -10 -36
rect -2 -38 2 -36
rect 10 -38 14 -36
<< ndiffusion >>
rect -17 -36 -14 -29
rect -10 -36 -9 -29
rect -4 -36 -2 -29
rect 2 -36 3 -29
rect 9 -36 10 -29
rect 14 -36 17 -29
rect 22 -36 26 -29
<< pdiffusion >>
rect -17 1 -14 8
rect -10 1 -2 8
rect 2 1 10 8
rect 14 1 17 8
rect 22 1 26 8
<< metal1 >>
rect -24 8 -17 20
rect -12 15 -7 20
rect -2 15 3 20
rect 8 15 11 20
rect 17 -12 22 1
rect -9 -17 22 -12
rect -9 -29 -4 -17
rect 17 -29 22 -17
rect -24 -46 -17 -36
rect 3 -41 9 -36
rect -12 -46 -7 -41
rect -2 -46 3 -41
rect 8 -46 11 -41
<< ntransistor >>
rect -14 -36 -10 -29
rect -2 -36 2 -29
rect 10 -36 14 -29
<< ptransistor >>
rect -14 1 -10 8
rect -2 1 2 8
rect 10 1 14 8
<< ndcontact >>
rect -24 -36 -17 -29
rect -9 -36 -4 -29
rect 3 -36 9 -29
rect 17 -36 22 -29
<< pdcontact >>
rect -24 1 -17 8
rect 17 1 22 8
<< psubstratepcontact >>
rect -17 -46 -12 -41
rect -7 -46 -2 -41
rect 3 -46 8 -41
<< nsubstratencontact >>
rect -17 15 -12 20
rect -7 15 -2 20
rect 3 15 8 20
<< labels >>
rlabel metal1 -21 17 -21 17 5 vdd!
rlabel metal1 -21 -43 -21 -43 1 gnd!
rlabel polysilicon -12 -3 -12 -3 1 a
rlabel polysilicon 0 -3 0 -3 1 b
rlabel polysilicon 12 -3 12 -3 1 c
rlabel metal1 20 -15 20 -15 1 out
<< end >>
