magic
tech scmos
timestamp 1596730447
<< nwell >>
rect -11 -1 15 16
<< polysilicon >>
rect -1 7 1 9
rect -1 -15 1 2
rect -1 -22 1 -19
<< ndiffusion >>
rect -2 -19 -1 -15
rect 1 -19 2 -15
<< pdiffusion >>
rect -3 2 -1 7
rect 1 2 2 7
<< metal1 >>
rect -11 11 -8 15
rect -4 11 0 15
rect 4 11 8 15
rect 12 11 15 15
rect -7 7 -3 11
rect 2 -6 6 2
rect -11 -10 -5 -6
rect 2 -10 15 -6
rect 2 -15 6 -10
rect -12 -29 -10 -25
rect -6 -29 -2 -19
rect 2 -29 6 -25
rect 10 -29 13 -25
<< ntransistor >>
rect -1 -19 1 -15
<< ptransistor >>
rect -1 2 1 7
<< polycontact >>
rect -5 -10 -1 -6
<< ndcontact >>
rect -6 -19 -2 -15
rect 2 -19 6 -15
<< pdcontact >>
rect -7 2 -3 7
rect 2 2 6 7
<< psubstratepcontact >>
rect -10 -29 -6 -25
rect -2 -29 2 -25
rect 6 -29 10 -25
<< nsubstratencontact >>
rect -8 11 -4 15
rect 0 11 4 15
rect 8 11 12 15
<< labels >>
rlabel metal1 13 13 13 13 6 vdd!
rlabel metal1 12 -27 12 -27 8 gnd!
rlabel metal1 -11 -10 -11 -6 3 in
rlabel metal1 15 -10 15 -6 7 out
<< end >>
